package JustBlinksNotTypeLevel_topEntity_types;


endpackage : JustBlinksNotTypeLevel_topEntity_types

